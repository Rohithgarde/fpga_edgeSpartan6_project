module upcnt(clk, rst);
